*hpddcc.sp
.subckt hpddcc y1 y2 y3 vbb x z	g='g' min='min'
.param L1='1*min'
.param L2='1*min'
.param L3='1*min'
.param L4='1*min'
.param L5='1*min'
.param L6='1*min'
.param L7='1*min'
.param L8='4*min'
.param L9='1*min'
.param L10='5*min'
.param L11='5*min'

.param W1='5*g'
.param W2='1*g'
.param W3='10*g'
.param W4='4*g'
.param W5='5*g'
.param W6='4*g'
.param W7='1*g'
.param W8='1*g'
.param W9='14*g'
.param W10='1*g'
.param W11='60*g'

*name	drain	gate	source	bulk	type dimension		source and drain area	  source and drain perimeter
m6n 	net1 	net1 	vdd 	vdd 	pfet L=L1 W='W1*L1' ad='W1*L1*5*L1' as='W1*L1*5*L1' pd='2*W1*L1+10*L1' ps='2*W1*L1+10*L1'
m7n 	net2 	net1 	vdd 	vdd 	pfet L=L1 W='W1*L1' ad='W1*L1*5*L1' as='W1*L1*5*L1' pd='2*W1*L1+10*L1' ps='2*W1*L1+10*L1'
m4p 	net7 	net8 	vdd 	vdd 	pfet L=L2 W='W2*L2' ad='W2*L2*5*L2' as='W2*L2*5*L2' pd='2*W2*L2+10*L2' ps='2*W2*L2+10*L2'
m5p 	net9 	net3 	vdd 	vdd 	pfet L=L2 W='W2*L2' ad='W2*L2*5*L2' as='W2*L2*5*L2' pd='2*W2*L2+10*L2' ps='2*W2*L2+10*L2'
m3p 	z 	net7 	net8 	vdd 	pfet L=L3 W='W3*L3' ad='W3*L3*5*L3' as='W3*L3*5*L3' pd='2*W3*L3+10*L3' ps='2*W3*L3+10*L3'
m2p 	net8 	net3 	vdd 	vdd 	pfet L=L3 W='W3*L3' ad='W3*L3*5*L3' as='W3*L3*5*L3' pd='2*W3*L3+10*L3' ps='2*W3*L3+10*L3'
m1p 	net3 	net3 	vdd 	vdd 	pfet L=L3 W='W3*L3' ad='W3*L3*5*L3' as='W3*L3*5*L3' pd='2*W3*L3+10*L3' ps='2*W3*L3+10*L3'
m8 	net5 	net12 	vdd 	vdd 	pfet L=L3 W='W3*L3' ad='W3*L3*5*L3' as='W3*L3*5*L3' pd='2*W3*L3+10*L3' ps='2*W3*L3+10*L3'
m13 	net10 	net13 	x 	vdd 	pfet L=L3 W='W3*L3' ad='W3*L3*5*L3' as='W3*L3*5*L3' pd='2*W3*L3+10*L3' ps='2*W3*L3+10*L3'
m12 	net13 	net13 	net6 	vdd 	pfet L=L3 W='W3*L3' ad='W3*L3*5*L3' as='W3*L3*5*L3' pd='2*W3*L3+10*L3' ps='2*W3*L3+10*L3'
m7 	net12 	net14 	vdd 	vdd 	pfet L=L4 W='W4*L4' ad='W4*L4*5*L4' as='W4*L4*5*L4' pd='2*W4*L4+10*L4' ps='2*W4*L4+10*L4'
m6 	net14 	net14 	vdd 	vdd 	pfet L=L4 W='W4*L4' ad='W4*L4*5*L4' as='W4*L4*5*L4' pd='2*W4*L4+10*L4' ps='2*W4*L4+10*L4'
m6p 	net9 	net9 	vss 	gnd 	nfet L=L5 W='W5*L5' ad='W5*L5*5*L5' as='W5*L5*5*L5' pd='2*W5*L5+10*L5' ps='2*W5*L5+10*L5'
m7p 	net7 	net9 	vss 	gnd 	nfet L=L5 W='W5*L5' ad='W5*L5*5*L5' as='W5*L5*5*L5' pd='2*W5*L5+10*L5' ps='2*W5*L5+10*L5'
m11 	net3 	net5 	x 	gnd 	nfet L=L6 W='W6*L6' ad='W6*L6*5*L6' as='W6*L6*5*L6' pd='2*W6*L6+10*L6' ps='2*W6*L6+10*L6'
m10 	net5 	net5 	net6 	gnd 	nfet L=L6 W='W6*L6' ad='W6*L6*5*L6' as='W6*L6*5*L6' pd='2*W6*L6+10*L6' ps='2*W6*L6+10*L6'
m3n 	z 	net2 	net11 	gnd 	nfet L=L6 W='W6*L6' ad='W6*L6*5*L6' as='W6*L6*5*L6' pd='2*W6*L6+10*L6' ps='2*W6*L6+10*L6'
m2n 	net11 	net10 	vss 	gnd 	nfet L=L6 W='W6*L6' ad='W6*L6*5*L6' as='W6*L6*5*L6' pd='2*W6*L6+10*L6' ps='2*W6*L6+10*L6'
m1n 	net10 	net10 	vss 	gnd 	nfet L=L6 W='W6*L6' ad='W6*L6*5*L6' as='W6*L6*5*L6' pd='2*W6*L6+10*L6' ps='2*W6*L6+10*L6'
m4n 	net2 	net11 	vss 	gnd 	nfet L=L7 W='W7*L7' ad='W7*L7*5*L7' as='W7*L7*5*L7' pd='2*W7*L7+10*L7' ps='2*W7*L7+10*L7'
m5n 	net1 	net10 	vss 	gnd 	nfet L=L7 W='W7*L7' ad='W7*L7*5*L7' as='W7*L7*5*L7' pd='2*W7*L7+10*L7' ps='2*W7*L7+10*L7'
m9 	net13 	vbb 	vss 	gnd 	nfet L=L8 W='W8*L8' ad='W8*L8*5*L8' as='W8*L8*5*L8' pd='2*W8*L8+10*L8' ps='2*W8*L8+10*L8'
m5d	net15 	vbb 	vss 	gnd 	nfet L=L9 W='W9*L9' ad='W9*L9*5*L9' as='W9*L9*5*L9' pd='2*W9*L9+10*L9' ps='2*W9*L9+10*L9'
m5c 	net16 	vbb 	vss 	gnd 	nfet L=L9 W='W9*L9' ad='W9*L9*5*L9' as='W9*L9*5*L9' pd='2*W9*L9+10*L9' ps='2*W9*L9+10*L9'
m5b 	net17 	vbb 	vss 	gnd 	nfet L=L9 W='W9*L9' ad='W9*L9*5*L9' as='W9*L9*5*L9' pd='2*W9*L9+10*L9' ps='2*W9*L9+10*L9'
m5a 	net18 	vbb 	vss 	gnd 	nfet L=L9 W='W9*L9' ad='W9*L9*5*L9' as='W9*L9*5*L9' pd='2*W9*L9+10*L9' ps='2*W9*L9+10*L9'
m4 	net12 	y1 	net15 	gnd 	nfet L=L10 W='W10*L10' ad='W10*L10*5*L10' as='W10*L10*5*L10' pd='2*W10*L10+10*L10' ps='2*W10*L10+10*L10'
m3 	net14 	x 	net16 	gnd 	nfet L=L10 W='W10*L10' ad='W10*L10*5*L10' as='W10*L10*5*L10' pd='2*W10*L10+10*L10' ps='2*W10*L10+10*L10'
m2 	net12 	y3 	net17 	gnd 	nfet L=L10 W='W10*L10' ad='W10*L10*5*L10' as='W10*L10*5*L10' pd='2*W10*L10+10*L10' ps='2*W10*L10+10*L10'
m1 	net14 	y2 	net18 	gnd 	nfet L=L10 W='W10*L10' ad='W10*L10*5*L10' as='W10*L10*5*L10' pd='2*W10*L10+10*L10' ps='2*W10*L10+10*L10'
m4a	vdd 	y1 	net16 	gnd 	nfet L=L11 W='W11*L11' ad='W11*L11*5*L11' as='W11*L11*5*L11' pd='2*W11*L11+10*L11' ps='2*W11*L11+10*L11'
m3a 	vdd 	x 	net15 	gnd 	nfet L=L11 W='W11*L11' ad='W11*L11*5*L11' as='W11*L11*5*L11' pd='2*W11*L11+10*L11' ps='2*W11*L11+10*L11'
m2a	vdd 	y3 	net18 	gnd 	nfet L=L11 W='W11*L11' ad='W11*L11*5*L11' as='W11*L11*5*L11' pd='2*W11*L11+10*L11' ps='2*W11*L11+10*L11'
m1a 	vdd 	y2 	net17 	gnd 	nfet L=L11 W='W11*L11' ad='W11*L11*5*L11' as='W11*L11*5*L11' pd='2*W11*L11+10*L11' ps='2*W11*L11+10*L11'
.ends
.end
