*test.sp
*----------------------------------------
*Parameters and models
*----------------------------------------
.include "~/cad/analog_computer/hspice/models/1.0u/models.sp"
.include "~/cad/analog_computer/hspice/models/0.5u/models.sp"
.include "~/cad/analog_computer/hspice/models/0.13u/model013.lib_inc"
.include "~/cad/analog_computer/hspice/models/0.09u/hspice_example.include_model"
.include "~/cad/analog_computer/hspice/models/0.05u/models.sp"

.end
